FourBitAdder